module Sopc(
  input   clock,
  input   reset
);
endmodule
