module Sopc(
  input   clock,
  input   reset,
  output  io_success
);
  assign io_success = 1'h0;
endmodule
